library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity find_track is
  port(
	  pos_row, pos_col : in  unsigned(9 downto 0);
		off_track        : out std_logic
  );
end find_track;

architecture synth of find_track is

begin
  off_track <= '1' when
		((pos_row = 10d"0" or pos_row = 10d"1") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"2" or pos_row = 10d"3") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"4" or pos_row = 10d"5") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"6" or pos_row = 10d"7") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"8" or pos_row = 10d"9") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"10" or pos_row = 10d"11") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"12" or pos_row = 10d"13") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"14" or pos_row = 10d"15") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"16" or pos_row = 10d"17") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"18" or pos_row = 10d"19") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"20" or pos_row = 10d"21") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"22" or pos_row = 10d"23") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"24" or pos_row = 10d"25") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"26" or pos_row = 10d"27") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"28" or pos_row = 10d"29") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"30" or pos_row = 10d"31") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"32" or pos_row = 10d"33") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"34" or pos_row = 10d"35") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"36" or pos_row = 10d"37") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"38" or pos_row = 10d"39") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"40" or pos_row = 10d"41") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"42" or pos_row = 10d"43") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"44" or pos_row = 10d"45") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"46" or pos_row = 10d"47") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"48" or pos_row = 10d"49") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"50" or pos_row = 10d"51") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"52" or pos_row = 10d"53") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"54" or pos_row = 10d"55") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"56" or pos_row = 10d"57") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"58" or pos_row = 10d"59") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"60" or pos_row = 10d"61") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"62" or pos_row = 10d"63") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"64" or pos_row = 10d"65") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"66" or pos_row = 10d"67") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"68" or pos_row = 10d"69") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"70" or pos_row = 10d"71") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"72" or pos_row = 10d"73") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"74" or pos_row = 10d"75") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"76" or pos_row = 10d"77") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"78" or pos_row = 10d"79") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"80" or pos_row = 10d"81") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"82" or pos_row = 10d"83") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"84" or pos_row = 10d"85") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"86" or pos_row = 10d"87") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"88" or pos_row = 10d"89") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"90" or pos_row = 10d"91") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"92" or pos_row = 10d"93") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"94" or pos_row = 10d"95") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"96" or pos_row = 10d"97") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"96" or pos_row = 10d"97") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"98" or pos_row = 10d"99") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"98" or pos_row = 10d"99") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"100" or pos_row = 10d"101") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"100" or pos_row = 10d"101") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"102" or pos_row = 10d"103") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"102" or pos_row = 10d"103") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"104" or pos_row = 10d"105") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"104" or pos_row = 10d"105") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"106" or pos_row = 10d"107") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"106" or pos_row = 10d"107") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"108" or pos_row = 10d"109") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"108" or pos_row = 10d"109") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"110" or pos_row = 10d"111") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"110" or pos_row = 10d"111") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"112" or pos_row = 10d"113") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"112" or pos_row = 10d"113") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"114" or pos_row = 10d"115") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"114" or pos_row = 10d"115") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"116" or pos_row = 10d"117") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"116" or pos_row = 10d"117") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"118" or pos_row = 10d"119") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"118" or pos_row = 10d"119") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"120" or pos_row = 10d"121") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"120" or pos_row = 10d"121") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"122" or pos_row = 10d"123") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"122" or pos_row = 10d"123") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"124" or pos_row = 10d"125") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"124" or pos_row = 10d"125") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"126" or pos_row = 10d"127") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"126" or pos_row = 10d"127") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"128" or pos_row = 10d"129") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"128" or pos_row = 10d"129") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"130" or pos_row = 10d"131") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"130" or pos_row = 10d"131") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"132" or pos_row = 10d"133") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"132" or pos_row = 10d"133") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"134" or pos_row = 10d"135") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"134" or pos_row = 10d"135") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"136" or pos_row = 10d"137") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"136" or pos_row = 10d"137") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"138" or pos_row = 10d"139") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"138" or pos_row = 10d"139") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"140" or pos_row = 10d"141") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"140" or pos_row = 10d"141") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"142" or pos_row = 10d"143") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"142" or pos_row = 10d"143") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"144" or pos_row = 10d"145") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"144" or pos_row = 10d"145") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"146" or pos_row = 10d"147") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"146" or pos_row = 10d"147") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"148" or pos_row = 10d"149") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"148" or pos_row = 10d"149") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"150" or pos_row = 10d"151") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"150" or pos_row = 10d"151") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"152" or pos_row = 10d"153") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"152" or pos_row = 10d"153") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"154" or pos_row = 10d"155") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"154" or pos_row = 10d"155") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"156" or pos_row = 10d"157") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"156" or pos_row = 10d"157") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"158" or pos_row = 10d"159") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"158" or pos_row = 10d"159") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"160" or pos_row = 10d"161") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"160" or pos_row = 10d"161") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"162" or pos_row = 10d"163") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"162" or pos_row = 10d"163") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"164" or pos_row = 10d"165") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"164" or pos_row = 10d"165") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"166" or pos_row = 10d"167") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"166" or pos_row = 10d"167") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"168" or pos_row = 10d"169") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"168" or pos_row = 10d"169") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"170" or pos_row = 10d"171") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"170" or pos_row = 10d"171") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"172" or pos_row = 10d"173") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"172" or pos_row = 10d"173") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"174" or pos_row = 10d"175") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"174" or pos_row = 10d"175") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"176" or pos_row = 10d"177") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"176" or pos_row = 10d"177") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"178" or pos_row = 10d"179") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"178" or pos_row = 10d"179") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"180" or pos_row = 10d"181") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"180" or pos_row = 10d"181") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"182" or pos_row = 10d"183") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"182" or pos_row = 10d"183") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"184" or pos_row = 10d"185") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"184" or pos_row = 10d"185") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"186" or pos_row = 10d"187") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"186" or pos_row = 10d"187") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"188" or pos_row = 10d"189") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"188" or pos_row = 10d"189") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"190" or pos_row = 10d"191") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"190" or pos_row = 10d"191") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"192" or pos_row = 10d"193") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"192" or pos_row = 10d"193") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"194" or pos_row = 10d"195") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"194" or pos_row = 10d"195") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"196" or pos_row = 10d"197") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"196" or pos_row = 10d"197") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"198" or pos_row = 10d"199") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"198" or pos_row = 10d"199") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"200" or pos_row = 10d"201") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"200" or pos_row = 10d"201") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"202" or pos_row = 10d"203") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"202" or pos_row = 10d"203") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"204" or pos_row = 10d"205") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"204" or pos_row = 10d"205") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"206" or pos_row = 10d"207") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"206" or pos_row = 10d"207") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"208" or pos_row = 10d"209") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"208" or pos_row = 10d"209") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"210" or pos_row = 10d"211") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"210" or pos_row = 10d"211") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"212" or pos_row = 10d"213") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"212" or pos_row = 10d"213") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"214" or pos_row = 10d"215") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"214" or pos_row = 10d"215") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"216" or pos_row = 10d"217") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"216" or pos_row = 10d"217") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"218" or pos_row = 10d"219") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"218" or pos_row = 10d"219") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"220" or pos_row = 10d"221") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"220" or pos_row = 10d"221") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"222" or pos_row = 10d"223") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"222" or pos_row = 10d"223") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"224" or pos_row = 10d"225") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"224" or pos_row = 10d"225") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"226" or pos_row = 10d"227") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"226" or pos_row = 10d"227") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"228" or pos_row = 10d"229") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"228" or pos_row = 10d"229") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"230" or pos_row = 10d"231") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"230" or pos_row = 10d"231") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"232" or pos_row = 10d"233") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"232" or pos_row = 10d"233") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"234" or pos_row = 10d"235") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"234" or pos_row = 10d"235") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"236" or pos_row = 10d"237") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"236" or pos_row = 10d"237") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"238" or pos_row = 10d"239") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"238" or pos_row = 10d"239") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"240" or pos_row = 10d"241") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"240" or pos_row = 10d"241") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"242" or pos_row = 10d"243") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"242" or pos_row = 10d"243") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"244" or pos_row = 10d"245") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"244" or pos_row = 10d"245") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"246" or pos_row = 10d"247") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"246" or pos_row = 10d"247") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"248" or pos_row = 10d"249") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"248" or pos_row = 10d"249") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"250" or pos_row = 10d"251") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"250" or pos_row = 10d"251") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"252" or pos_row = 10d"253") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"252" or pos_row = 10d"253") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"254" or pos_row = 10d"255") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"254" or pos_row = 10d"255") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"256" or pos_row = 10d"257") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"256" or pos_row = 10d"257") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"258" or pos_row = 10d"259") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"258" or pos_row = 10d"259") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"260" or pos_row = 10d"261") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"260" or pos_row = 10d"261") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"262" or pos_row = 10d"263") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"262" or pos_row = 10d"263") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"264" or pos_row = 10d"265") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"264" or pos_row = 10d"265") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"266" or pos_row = 10d"267") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"266" or pos_row = 10d"267") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"268" or pos_row = 10d"269") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"268" or pos_row = 10d"269") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"270" or pos_row = 10d"271") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"270" or pos_row = 10d"271") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"272" or pos_row = 10d"273") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"272" or pos_row = 10d"273") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"274" or pos_row = 10d"275") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"274" or pos_row = 10d"275") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"276" or pos_row = 10d"277") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"276" or pos_row = 10d"277") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"278" or pos_row = 10d"279") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"278" or pos_row = 10d"279") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"280" or pos_row = 10d"281") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"280" or pos_row = 10d"281") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"282" or pos_row = 10d"283") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"282" or pos_row = 10d"283") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"284" or pos_row = 10d"285") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"284" or pos_row = 10d"285") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"286" or pos_row = 10d"287") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"286" or pos_row = 10d"287") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"288" or pos_row = 10d"289") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"288" or pos_row = 10d"289") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"290" or pos_row = 10d"291") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"290" or pos_row = 10d"291") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"292" or pos_row = 10d"293") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"292" or pos_row = 10d"293") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"294" or pos_row = 10d"295") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"294" or pos_row = 10d"295") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"296" or pos_row = 10d"297") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"296" or pos_row = 10d"297") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"298" or pos_row = 10d"299") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"298" or pos_row = 10d"299") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"300" or pos_row = 10d"301") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"300" or pos_row = 10d"301") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"302" or pos_row = 10d"303") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"302" or pos_row = 10d"303") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"304" or pos_row = 10d"305") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"304" or pos_row = 10d"305") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"306" or pos_row = 10d"307") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"306" or pos_row = 10d"307") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"308" or pos_row = 10d"309") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"308" or pos_row = 10d"309") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"310" or pos_row = 10d"311") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"310" or pos_row = 10d"311") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"312" or pos_row = 10d"313") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"312" or pos_row = 10d"313") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"314" or pos_row = 10d"315") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"314" or pos_row = 10d"315") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"316" or pos_row = 10d"317") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"316" or pos_row = 10d"317") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"318" or pos_row = 10d"319") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"318" or pos_row = 10d"319") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"320" or pos_row = 10d"321") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"320" or pos_row = 10d"321") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"322" or pos_row = 10d"323") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"322" or pos_row = 10d"323") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"324" or pos_row = 10d"325") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"324" or pos_row = 10d"325") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"326" or pos_row = 10d"327") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"326" or pos_row = 10d"327") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"328" or pos_row = 10d"329") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"328" or pos_row = 10d"329") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"330" or pos_row = 10d"331") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"330" or pos_row = 10d"331") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"332" or pos_row = 10d"333") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"332" or pos_row = 10d"333") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"334" or pos_row = 10d"335") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"334" or pos_row = 10d"335") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"336" or pos_row = 10d"337") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"336" or pos_row = 10d"337") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"338" or pos_row = 10d"339") and (pos_col >= 10d"0" and pos_col < 10d"150")) or
		((pos_row = 10d"338" or pos_row = 10d"339") and (pos_col >= 10d"500" and pos_col < 10d"640")) or
		((pos_row = 10d"340" or pos_row = 10d"341") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"342" or pos_row = 10d"343") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"344" or pos_row = 10d"345") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"346" or pos_row = 10d"347") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"348" or pos_row = 10d"349") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"350" or pos_row = 10d"351") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"352" or pos_row = 10d"353") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"354" or pos_row = 10d"355") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"356" or pos_row = 10d"357") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"358" or pos_row = 10d"359") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"360" or pos_row = 10d"361") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"362" or pos_row = 10d"363") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"364" or pos_row = 10d"365") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"366" or pos_row = 10d"367") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"368" or pos_row = 10d"369") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"370" or pos_row = 10d"371") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"372" or pos_row = 10d"373") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"374" or pos_row = 10d"375") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"376" or pos_row = 10d"377") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"378" or pos_row = 10d"379") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"380" or pos_row = 10d"381") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"382" or pos_row = 10d"383") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"384" or pos_row = 10d"385") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"386" or pos_row = 10d"387") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"388" or pos_row = 10d"389") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"390" or pos_row = 10d"391") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"392" or pos_row = 10d"393") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"394" or pos_row = 10d"395") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"396" or pos_row = 10d"397") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"398" or pos_row = 10d"399") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"400" or pos_row = 10d"401") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"402" or pos_row = 10d"403") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"404" or pos_row = 10d"405") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"406" or pos_row = 10d"407") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"408" or pos_row = 10d"409") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"410" or pos_row = 10d"411") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"412" or pos_row = 10d"413") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"414" or pos_row = 10d"415") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"416" or pos_row = 10d"417") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"418" or pos_row = 10d"419") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"420" or pos_row = 10d"421") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"422" or pos_row = 10d"423") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"424" or pos_row = 10d"425") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"426" or pos_row = 10d"427") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"428" or pos_row = 10d"429") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"430" or pos_row = 10d"431") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"432" or pos_row = 10d"433") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"434" or pos_row = 10d"435") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"436" or pos_row = 10d"437") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"438" or pos_row = 10d"439") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"440" or pos_row = 10d"441") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"442" or pos_row = 10d"443") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"444" or pos_row = 10d"445") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"446" or pos_row = 10d"447") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"448" or pos_row = 10d"449") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"450" or pos_row = 10d"451") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"452" or pos_row = 10d"453") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"454" or pos_row = 10d"455") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"456" or pos_row = 10d"457") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"458" or pos_row = 10d"459") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"460" or pos_row = 10d"461") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"462" or pos_row = 10d"463") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"464" or pos_row = 10d"465") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"466" or pos_row = 10d"467") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"468" or pos_row = 10d"469") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"470" or pos_row = 10d"471") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"472" or pos_row = 10d"473") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"474" or pos_row = 10d"475") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"476" or pos_row = 10d"477") and (pos_col >= 10d"0" and pos_col < 10d"640")) or
		((pos_row = 10d"478" or pos_row = 10d"479") and (pos_col >= 10d"0" and pos_col < 10d"640")) else '0';
end;
