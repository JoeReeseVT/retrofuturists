library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity win_rgb is
  port(
		player	: in std_logic;
    vga_row : in  unsigned(9 downto 0);
		vga_col : in  unsigned(9 downto 0);
		
    rgb_o   : out std_logic_vector(5 downto 0)
  );
end win_rgb;

architecture synth of win_rgb is

begin

rgb_o <= "110000" when player = '0' and 
								(((vga_row >= 10d"152" and vga_row < 10d"156") and (vga_col >= 10d"124" and vga_col < 10d"136")) or
								((vga_row >= 10d"152" and vga_row < 10d"156") and (vga_col >= 10d"160" and vga_col < 10d"172")) or
								((vga_row >= 10d"152" and vga_row < 10d"156") and (vga_col >= 10d"196" and vga_col < 10d"208")) or
								((vga_row >= 10d"152" and vga_row < 10d"156") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"152" and vga_row < 10d"156") and (vga_col >= 10d"236" and vga_col < 10d"248")) or
								((vga_row >= 10d"152" and vga_row < 10d"156") and (vga_col >= 10d"276" and vga_col < 10d"288")) or
								((vga_row >= 10d"152" and vga_row < 10d"156") and (vga_col >= 10d"304" and vga_col < 10d"316")) or
								((vga_row >= 10d"152" and vga_row < 10d"156") and (vga_col >= 10d"344" and vga_col < 10d"356")) or
								((vga_row >= 10d"152" and vga_row < 10d"156") and (vga_col >= 10d"372" and vga_col < 10d"420")) or
								((vga_row >= 10d"152" and vga_row < 10d"156") and (vga_col >= 10d"432" and vga_col < 10d"476")) or
								((vga_row >= 10d"156" and vga_row < 10d"160") and (vga_col >= 10d"124" and vga_col < 10d"136")) or
								((vga_row >= 10d"156" and vga_row < 10d"160") and (vga_col >= 10d"160" and vga_col < 10d"172")) or
								((vga_row >= 10d"156" and vga_row < 10d"160") and (vga_col >= 10d"196" and vga_col < 10d"208")) or
								((vga_row >= 10d"156" and vga_row < 10d"160") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"156" and vga_row < 10d"160") and (vga_col >= 10d"236" and vga_col < 10d"252")) or
								((vga_row >= 10d"156" and vga_row < 10d"160") and (vga_col >= 10d"276" and vga_col < 10d"288")) or
								((vga_row >= 10d"156" and vga_row < 10d"160") and (vga_col >= 10d"304" and vga_col < 10d"320")) or
								((vga_row >= 10d"156" and vga_row < 10d"160") and (vga_col >= 10d"344" and vga_col < 10d"356")) or
								((vga_row >= 10d"156" and vga_row < 10d"160") and (vga_col >= 10d"372" and vga_col < 10d"420")) or
								((vga_row >= 10d"156" and vga_row < 10d"160") and (vga_col >= 10d"432" and vga_col < 10d"480")) or
								((vga_row >= 10d"160" and vga_row < 10d"164") and (vga_col >= 10d"128" and vga_col < 10d"140")) or
								((vga_row >= 10d"160" and vga_row < 10d"164") and (vga_col >= 10d"156" and vga_col < 10d"176")) or
								((vga_row >= 10d"160" and vga_row < 10d"164") and (vga_col >= 10d"192" and vga_col < 10d"204")) or
								((vga_row >= 10d"160" and vga_row < 10d"164") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"160" and vga_row < 10d"164") and (vga_col >= 10d"236" and vga_col < 10d"256")) or
								((vga_row >= 10d"160" and vga_row < 10d"164") and (vga_col >= 10d"276" and vga_col < 10d"288")) or
								((vga_row >= 10d"160" and vga_row < 10d"164") and (vga_col >= 10d"304" and vga_col < 10d"324")) or
								((vga_row >= 10d"160" and vga_row < 10d"164") and (vga_col >= 10d"344" and vga_col < 10d"356")) or
								((vga_row >= 10d"160" and vga_row < 10d"164") and (vga_col >= 10d"372" and vga_col < 10d"420")) or
								((vga_row >= 10d"160" and vga_row < 10d"164") and (vga_col >= 10d"432" and vga_col < 10d"484")) or
								((vga_row >= 10d"164" and vga_row < 10d"168") and (vga_col >= 10d"128" and vga_col < 10d"140")) or
								((vga_row >= 10d"164" and vga_row < 10d"168") and (vga_col >= 10d"156" and vga_col < 10d"176")) or
								((vga_row >= 10d"164" and vga_row < 10d"168") and (vga_col >= 10d"192" and vga_col < 10d"204")) or
								((vga_row >= 10d"164" and vga_row < 10d"168") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"164" and vga_row < 10d"168") and (vga_col >= 10d"236" and vga_col < 10d"256")) or
								((vga_row >= 10d"164" and vga_row < 10d"168") and (vga_col >= 10d"276" and vga_col < 10d"288")) or
								((vga_row >= 10d"164" and vga_row < 10d"168") and (vga_col >= 10d"304" and vga_col < 10d"324")) or
								((vga_row >= 10d"164" and vga_row < 10d"168") and (vga_col >= 10d"344" and vga_col < 10d"356")) or
								((vga_row >= 10d"164" and vga_row < 10d"168") and (vga_col >= 10d"372" and vga_col < 10d"384")) or
								((vga_row >= 10d"164" and vga_row < 10d"168") and (vga_col >= 10d"432" and vga_col < 10d"444")) or
								((vga_row >= 10d"164" and vga_row < 10d"168") and (vga_col >= 10d"468" and vga_col < 10d"484")) or
								((vga_row >= 10d"168" and vga_row < 10d"172") and (vga_col >= 10d"128" and vga_col < 10d"140")) or
								((vga_row >= 10d"168" and vga_row < 10d"172") and (vga_col >= 10d"156" and vga_col < 10d"164")) or
								((vga_row >= 10d"168" and vga_row < 10d"172") and (vga_col >= 10d"168" and vga_col < 10d"176")) or
								((vga_row >= 10d"168" and vga_row < 10d"172") and (vga_col >= 10d"192" and vga_col < 10d"204")) or
								((vga_row >= 10d"168" and vga_row < 10d"172") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"168" and vga_row < 10d"172") and (vga_col >= 10d"236" and vga_col < 10d"260")) or
								((vga_row >= 10d"168" and vga_row < 10d"172") and (vga_col >= 10d"276" and vga_col < 10d"288")) or
								((vga_row >= 10d"168" and vga_row < 10d"172") and (vga_col >= 10d"304" and vga_col < 10d"328")) or
								((vga_row >= 10d"168" and vga_row < 10d"172") and (vga_col >= 10d"344" and vga_col < 10d"356")) or
								((vga_row >= 10d"168" and vga_row < 10d"172") and (vga_col >= 10d"372" and vga_col < 10d"384")) or
								((vga_row >= 10d"168" and vga_row < 10d"172") and (vga_col >= 10d"432" and vga_col < 10d"444")) or
								((vga_row >= 10d"168" and vga_row < 10d"172") and (vga_col >= 10d"472" and vga_col < 10d"484")) or
								((vga_row >= 10d"172" and vga_row < 10d"176") and (vga_col >= 10d"128" and vga_col < 10d"140")) or
								((vga_row >= 10d"172" and vga_row < 10d"176") and (vga_col >= 10d"152" and vga_col < 10d"164")) or
								((vga_row >= 10d"172" and vga_row < 10d"176") and (vga_col >= 10d"168" and vga_col < 10d"180")) or
								((vga_row >= 10d"172" and vga_row < 10d"176") and (vga_col >= 10d"192" and vga_col < 10d"204")) or
								((vga_row >= 10d"172" and vga_row < 10d"176") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"172" and vga_row < 10d"176") and (vga_col >= 10d"236" and vga_col < 10d"260")) or
								((vga_row >= 10d"172" and vga_row < 10d"176") and (vga_col >= 10d"276" and vga_col < 10d"288")) or
								((vga_row >= 10d"172" and vga_row < 10d"176") and (vga_col >= 10d"304" and vga_col < 10d"328")) or
								((vga_row >= 10d"172" and vga_row < 10d"176") and (vga_col >= 10d"344" and vga_col < 10d"356")) or
								((vga_row >= 10d"172" and vga_row < 10d"176") and (vga_col >= 10d"372" and vga_col < 10d"384")) or
								((vga_row >= 10d"172" and vga_row < 10d"176") and (vga_col >= 10d"432" and vga_col < 10d"444")) or
								((vga_row >= 10d"172" and vga_row < 10d"176") and (vga_col >= 10d"472" and vga_col < 10d"484")) or
								((vga_row >= 10d"172" and vga_row < 10d"176") and (vga_col >= 10d"500" and vga_col < 10d"512")) or
								((vga_row >= 10d"176" and vga_row < 10d"180") and (vga_col >= 10d"128" and vga_col < 10d"140")) or
								((vga_row >= 10d"176" and vga_row < 10d"180") and (vga_col >= 10d"152" and vga_col < 10d"164")) or
								((vga_row >= 10d"176" and vga_row < 10d"180") and (vga_col >= 10d"168" and vga_col < 10d"180")) or
								((vga_row >= 10d"176" and vga_row < 10d"180") and (vga_col >= 10d"192" and vga_col < 10d"204")) or
								((vga_row >= 10d"176" and vga_row < 10d"180") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"176" and vga_row < 10d"180") and (vga_col >= 10d"236" and vga_col < 10d"248")) or
								((vga_row >= 10d"176" and vga_row < 10d"180") and (vga_col >= 10d"252" and vga_col < 10d"264")) or
								((vga_row >= 10d"176" and vga_row < 10d"180") and (vga_col >= 10d"276" and vga_col < 10d"288")) or
								((vga_row >= 10d"176" and vga_row < 10d"180") and (vga_col >= 10d"304" and vga_col < 10d"316")) or
								((vga_row >= 10d"176" and vga_row < 10d"180") and (vga_col >= 10d"320" and vga_col < 10d"332")) or
								((vga_row >= 10d"176" and vga_row < 10d"180") and (vga_col >= 10d"344" and vga_col < 10d"356")) or
								((vga_row >= 10d"176" and vga_row < 10d"180") and (vga_col >= 10d"372" and vga_col < 10d"384")) or
								((vga_row >= 10d"176" and vga_row < 10d"180") and (vga_col >= 10d"432" and vga_col < 10d"444")) or
								((vga_row >= 10d"176" and vga_row < 10d"180") and (vga_col >= 10d"468" and vga_col < 10d"484")) or
								((vga_row >= 10d"176" and vga_row < 10d"180") and (vga_col >= 10d"500" and vga_col < 10d"512")) or
								((vga_row >= 10d"180" and vga_row < 10d"184") and (vga_col >= 10d"132" and vga_col < 10d"144")) or
								((vga_row >= 10d"180" and vga_row < 10d"184") and (vga_col >= 10d"152" and vga_col < 10d"164")) or
								((vga_row >= 10d"180" and vga_row < 10d"184") and (vga_col >= 10d"168" and vga_col < 10d"180")) or
								((vga_row >= 10d"180" and vga_row < 10d"184") and (vga_col >= 10d"188" and vga_col < 10d"200")) or
								((vga_row >= 10d"180" and vga_row < 10d"184") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"180" and vga_row < 10d"184") and (vga_col >= 10d"236" and vga_col < 10d"248")) or
								((vga_row >= 10d"180" and vga_row < 10d"184") and (vga_col >= 10d"252" and vga_col < 10d"264")) or
								((vga_row >= 10d"180" and vga_row < 10d"184") and (vga_col >= 10d"276" and vga_col < 10d"288")) or
								((vga_row >= 10d"180" and vga_row < 10d"184") and (vga_col >= 10d"304" and vga_col < 10d"316")) or
								((vga_row >= 10d"180" and vga_row < 10d"184") and (vga_col >= 10d"320" and vga_col < 10d"332")) or
								((vga_row >= 10d"180" and vga_row < 10d"184") and (vga_col >= 10d"344" and vga_col < 10d"356")) or
								((vga_row >= 10d"180" and vga_row < 10d"184") and (vga_col >= 10d"372" and vga_col < 10d"416")) or
								((vga_row >= 10d"180" and vga_row < 10d"184") and (vga_col >= 10d"432" and vga_col < 10d"480")) or
								((vga_row >= 10d"180" and vga_row < 10d"184") and (vga_col >= 10d"500" and vga_col < 10d"512")) or
								((vga_row >= 10d"184" and vga_row < 10d"188") and (vga_col >= 10d"132" and vga_col < 10d"144")) or
								((vga_row >= 10d"184" and vga_row < 10d"188") and (vga_col >= 10d"148" and vga_col < 10d"160")) or
								((vga_row >= 10d"184" and vga_row < 10d"188") and (vga_col >= 10d"172" and vga_col < 10d"180")) or
								((vga_row >= 10d"184" and vga_row < 10d"188") and (vga_col >= 10d"188" and vga_col < 10d"200")) or
								((vga_row >= 10d"184" and vga_row < 10d"188") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"184" and vga_row < 10d"188") and (vga_col >= 10d"236" and vga_col < 10d"248")) or
								((vga_row >= 10d"184" and vga_row < 10d"188") and (vga_col >= 10d"256" and vga_col < 10d"268")) or
								((vga_row >= 10d"184" and vga_row < 10d"188") and (vga_col >= 10d"276" and vga_col < 10d"288")) or
								((vga_row >= 10d"184" and vga_row < 10d"188") and (vga_col >= 10d"304" and vga_col < 10d"316")) or
								((vga_row >= 10d"184" and vga_row < 10d"188") and (vga_col >= 10d"324" and vga_col < 10d"336")) or
								((vga_row >= 10d"184" and vga_row < 10d"188") and (vga_col >= 10d"344" and vga_col < 10d"356")) or
								((vga_row >= 10d"184" and vga_row < 10d"188") and (vga_col >= 10d"372" and vga_col < 10d"416")) or
								((vga_row >= 10d"184" and vga_row < 10d"188") and (vga_col >= 10d"432" and vga_col < 10d"476")) or
								((vga_row >= 10d"188" and vga_row < 10d"192") and (vga_col >= 10d"132" and vga_col < 10d"144")) or
								((vga_row >= 10d"188" and vga_row < 10d"192") and (vga_col >= 10d"148" and vga_col < 10d"160")) or
								((vga_row >= 10d"188" and vga_row < 10d"192") and (vga_col >= 10d"172" and vga_col < 10d"184")) or
								((vga_row >= 10d"188" and vga_row < 10d"192") and (vga_col >= 10d"188" and vga_col < 10d"200")) or
								((vga_row >= 10d"188" and vga_row < 10d"192") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"188" and vga_row < 10d"192") and (vga_col >= 10d"236" and vga_col < 10d"248")) or
								((vga_row >= 10d"188" and vga_row < 10d"192") and (vga_col >= 10d"256" and vga_col < 10d"272")) or
								((vga_row >= 10d"188" and vga_row < 10d"192") and (vga_col >= 10d"276" and vga_col < 10d"288")) or
								((vga_row >= 10d"188" and vga_row < 10d"192") and (vga_col >= 10d"304" and vga_col < 10d"316")) or
								((vga_row >= 10d"188" and vga_row < 10d"192") and (vga_col >= 10d"324" and vga_col < 10d"340")) or
								((vga_row >= 10d"188" and vga_row < 10d"192") and (vga_col >= 10d"344" and vga_col < 10d"356")) or
								((vga_row >= 10d"188" and vga_row < 10d"192") and (vga_col >= 10d"372" and vga_col < 10d"416")) or
								((vga_row >= 10d"188" and vga_row < 10d"192") and (vga_col >= 10d"432" and vga_col < 10d"468")) or
								((vga_row >= 10d"192" and vga_row < 10d"196") and (vga_col >= 10d"132" and vga_col < 10d"144")) or
								((vga_row >= 10d"192" and vga_row < 10d"196") and (vga_col >= 10d"148" and vga_col < 10d"160")) or
								((vga_row >= 10d"192" and vga_row < 10d"196") and (vga_col >= 10d"172" and vga_col < 10d"184")) or
								((vga_row >= 10d"192" and vga_row < 10d"196") and (vga_col >= 10d"188" and vga_col < 10d"200")) or
								((vga_row >= 10d"192" and vga_row < 10d"196") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"192" and vga_row < 10d"196") and (vga_col >= 10d"236" and vga_col < 10d"248")) or
								((vga_row >= 10d"192" and vga_row < 10d"196") and (vga_col >= 10d"260" and vga_col < 10d"272")) or
								((vga_row >= 10d"192" and vga_row < 10d"196") and (vga_col >= 10d"276" and vga_col < 10d"288")) or
								((vga_row >= 10d"192" and vga_row < 10d"196") and (vga_col >= 10d"304" and vga_col < 10d"316")) or
								((vga_row >= 10d"192" and vga_row < 10d"196") and (vga_col >= 10d"328" and vga_col < 10d"340")) or
								((vga_row >= 10d"192" and vga_row < 10d"196") and (vga_col >= 10d"344" and vga_col < 10d"356")) or
								((vga_row >= 10d"192" and vga_row < 10d"196") and (vga_col >= 10d"372" and vga_col < 10d"384")) or
								((vga_row >= 10d"192" and vga_row < 10d"196") and (vga_col >= 10d"432" and vga_col < 10d"444")) or
								((vga_row >= 10d"192" and vga_row < 10d"196") and (vga_col >= 10d"456" and vga_col < 10d"472")) or
								((vga_row >= 10d"196" and vga_row < 10d"200") and (vga_col >= 10d"136" and vga_col < 10d"144")) or
								((vga_row >= 10d"196" and vga_row < 10d"200") and (vga_col >= 10d"148" and vga_col < 10d"160")) or
								((vga_row >= 10d"196" and vga_row < 10d"200") and (vga_col >= 10d"172" and vga_col < 10d"184")) or
								((vga_row >= 10d"196" and vga_row < 10d"200") and (vga_col >= 10d"188" and vga_col < 10d"196")) or
								((vga_row >= 10d"196" and vga_row < 10d"200") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"196" and vga_row < 10d"200") and (vga_col >= 10d"236" and vga_col < 10d"248")) or
								((vga_row >= 10d"196" and vga_row < 10d"200") and (vga_col >= 10d"264" and vga_col < 10d"288")) or
								((vga_row >= 10d"196" and vga_row < 10d"200") and (vga_col >= 10d"304" and vga_col < 10d"316")) or
								((vga_row >= 10d"196" and vga_row < 10d"200") and (vga_col >= 10d"332" and vga_col < 10d"356")) or
								((vga_row >= 10d"196" and vga_row < 10d"200") and (vga_col >= 10d"372" and vga_col < 10d"384")) or
								((vga_row >= 10d"196" and vga_row < 10d"200") and (vga_col >= 10d"432" and vga_col < 10d"444")) or
								((vga_row >= 10d"196" and vga_row < 10d"200") and (vga_col >= 10d"460" and vga_col < 10d"476")) or
								((vga_row >= 10d"200" and vga_row < 10d"204") and (vga_col >= 10d"136" and vga_col < 10d"156")) or
								((vga_row >= 10d"200" and vga_row < 10d"204") and (vga_col >= 10d"176" and vga_col < 10d"196")) or
								((vga_row >= 10d"200" and vga_row < 10d"204") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"200" and vga_row < 10d"204") and (vga_col >= 10d"236" and vga_col < 10d"248")) or
								((vga_row >= 10d"200" and vga_row < 10d"204") and (vga_col >= 10d"264" and vga_col < 10d"288")) or
								((vga_row >= 10d"200" and vga_row < 10d"204") and (vga_col >= 10d"304" and vga_col < 10d"316")) or
								((vga_row >= 10d"200" and vga_row < 10d"204") and (vga_col >= 10d"332" and vga_col < 10d"356")) or
								((vga_row >= 10d"200" and vga_row < 10d"204") and (vga_col >= 10d"372" and vga_col < 10d"384")) or
								((vga_row >= 10d"200" and vga_row < 10d"204") and (vga_col >= 10d"432" and vga_col < 10d"444")) or
								((vga_row >= 10d"200" and vga_row < 10d"204") and (vga_col >= 10d"464" and vga_col < 10d"476")) or
								((vga_row >= 10d"204" and vga_row < 10d"208") and (vga_col >= 10d"136" and vga_col < 10d"156")) or
								((vga_row >= 10d"204" and vga_row < 10d"208") and (vga_col >= 10d"176" and vga_col < 10d"196")) or
								((vga_row >= 10d"204" and vga_row < 10d"208") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"204" and vga_row < 10d"208") and (vga_col >= 10d"236" and vga_col < 10d"248")) or
								((vga_row >= 10d"204" and vga_row < 10d"208") and (vga_col >= 10d"268" and vga_col < 10d"288")) or
								((vga_row >= 10d"204" and vga_row < 10d"208") and (vga_col >= 10d"304" and vga_col < 10d"316")) or
								((vga_row >= 10d"204" and vga_row < 10d"208") and (vga_col >= 10d"336" and vga_col < 10d"356")) or
								((vga_row >= 10d"204" and vga_row < 10d"208") and (vga_col >= 10d"372" and vga_col < 10d"384")) or
								((vga_row >= 10d"204" and vga_row < 10d"208") and (vga_col >= 10d"432" and vga_col < 10d"444")) or
								((vga_row >= 10d"204" and vga_row < 10d"208") and (vga_col >= 10d"468" and vga_col < 10d"480")) or
								((vga_row >= 10d"208" and vga_row < 10d"212") and (vga_col >= 10d"136" and vga_col < 10d"156")) or
								((vga_row >= 10d"208" and vga_row < 10d"212") and (vga_col >= 10d"176" and vga_col < 10d"196")) or
								((vga_row >= 10d"208" and vga_row < 10d"212") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"208" and vga_row < 10d"212") and (vga_col >= 10d"236" and vga_col < 10d"248")) or
								((vga_row >= 10d"208" and vga_row < 10d"212") and (vga_col >= 10d"268" and vga_col < 10d"288")) or
								((vga_row >= 10d"208" and vga_row < 10d"212") and (vga_col >= 10d"304" and vga_col < 10d"316")) or
								((vga_row >= 10d"208" and vga_row < 10d"212") and (vga_col >= 10d"336" and vga_col < 10d"356")) or
								((vga_row >= 10d"208" and vga_row < 10d"212") and (vga_col >= 10d"372" and vga_col < 10d"420")) or
								((vga_row >= 10d"208" and vga_row < 10d"212") and (vga_col >= 10d"432" and vga_col < 10d"444")) or
								((vga_row >= 10d"208" and vga_row < 10d"212") and (vga_col >= 10d"468" and vga_col < 10d"484")) or
								((vga_row >= 10d"208" and vga_row < 10d"212") and (vga_col >= 10d"500" and vga_col < 10d"512")) or
								((vga_row >= 10d"212" and vga_row < 10d"216") and (vga_col >= 10d"140" and vga_col < 10d"152")) or
								((vga_row >= 10d"212" and vga_row < 10d"216") and (vga_col >= 10d"180" and vga_col < 10d"192")) or
								((vga_row >= 10d"212" and vga_row < 10d"216") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"212" and vga_row < 10d"216") and (vga_col >= 10d"236" and vga_col < 10d"248")) or
								((vga_row >= 10d"212" and vga_row < 10d"216") and (vga_col >= 10d"272" and vga_col < 10d"288")) or
								((vga_row >= 10d"212" and vga_row < 10d"216") and (vga_col >= 10d"304" and vga_col < 10d"316")) or
								((vga_row >= 10d"212" and vga_row < 10d"216") and (vga_col >= 10d"340" and vga_col < 10d"356")) or
								((vga_row >= 10d"212" and vga_row < 10d"216") and (vga_col >= 10d"372" and vga_col < 10d"420")) or
								((vga_row >= 10d"212" and vga_row < 10d"216") and (vga_col >= 10d"432" and vga_col < 10d"444")) or
								((vga_row >= 10d"212" and vga_row < 10d"216") and (vga_col >= 10d"472" and vga_col < 10d"484")) or
								((vga_row >= 10d"212" and vga_row < 10d"216") and (vga_col >= 10d"500" and vga_col < 10d"512")) or
								((vga_row >= 10d"216" and vga_row < 10d"220") and (vga_col >= 10d"140" and vga_col < 10d"152")) or
								((vga_row >= 10d"216" and vga_row < 10d"220") and (vga_col >= 10d"180" and vga_col < 10d"192")) or
								((vga_row >= 10d"216" and vga_row < 10d"220") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"216" and vga_row < 10d"220") and (vga_col >= 10d"236" and vga_col < 10d"248")) or
								((vga_row >= 10d"216" and vga_row < 10d"220") and (vga_col >= 10d"272" and vga_col < 10d"288")) or
								((vga_row >= 10d"216" and vga_row < 10d"220") and (vga_col >= 10d"304" and vga_col < 10d"316")) or
								((vga_row >= 10d"216" and vga_row < 10d"220") and (vga_col >= 10d"340" and vga_col < 10d"356")) or
								((vga_row >= 10d"216" and vga_row < 10d"220") and (vga_col >= 10d"372" and vga_col < 10d"420")) or
								((vga_row >= 10d"216" and vga_row < 10d"220") and (vga_col >= 10d"432" and vga_col < 10d"444")) or
								((vga_row >= 10d"216" and vga_row < 10d"220") and (vga_col >= 10d"472" and vga_col < 10d"488")) or
								((vga_row >= 10d"216" and vga_row < 10d"220") and (vga_col >= 10d"500" and vga_col < 10d"512")) or
								((vga_row >= 10d"256" and vga_row < 10d"260") and (vga_col >= 10d"232" and vga_col < 10d"276")) or
								((vga_row >= 10d"256" and vga_row < 10d"260") and (vga_col >= 10d"300" and vga_col < 10d"348")) or
								((vga_row >= 10d"256" and vga_row < 10d"260") and (vga_col >= 10d"360" and vga_col < 10d"400")) or
								((vga_row >= 10d"260" and vga_row < 10d"264") and (vga_col >= 10d"232" and vga_col < 10d"280")) or
								((vga_row >= 10d"260" and vga_row < 10d"264") and (vga_col >= 10d"300" and vga_col < 10d"348")) or
								((vga_row >= 10d"260" and vga_row < 10d"264") and (vga_col >= 10d"360" and vga_col < 10d"404")) or
								((vga_row >= 10d"264" and vga_row < 10d"268") and (vga_col >= 10d"232" and vga_col < 10d"284")) or
								((vga_row >= 10d"264" and vga_row < 10d"268") and (vga_col >= 10d"300" and vga_col < 10d"348")) or
								((vga_row >= 10d"264" and vga_row < 10d"268") and (vga_col >= 10d"360" and vga_col < 10d"408")) or
								((vga_row >= 10d"268" and vga_row < 10d"272") and (vga_col >= 10d"232" and vga_col < 10d"244")) or
								((vga_row >= 10d"268" and vga_row < 10d"272") and (vga_col >= 10d"268" and vga_col < 10d"284")) or
								((vga_row >= 10d"268" and vga_row < 10d"272") and (vga_col >= 10d"300" and vga_col < 10d"312")) or
								((vga_row >= 10d"268" and vga_row < 10d"272") and (vga_col >= 10d"360" and vga_col < 10d"372")) or
								((vga_row >= 10d"268" and vga_row < 10d"272") and (vga_col >= 10d"396" and vga_col < 10d"412")) or
								((vga_row >= 10d"272" and vga_row < 10d"276") and (vga_col >= 10d"232" and vga_col < 10d"244")) or
								((vga_row >= 10d"272" and vga_row < 10d"276") and (vga_col >= 10d"272" and vga_col < 10d"284")) or
								((vga_row >= 10d"272" and vga_row < 10d"276") and (vga_col >= 10d"300" and vga_col < 10d"312")) or
								((vga_row >= 10d"272" and vga_row < 10d"276") and (vga_col >= 10d"360" and vga_col < 10d"372")) or
								((vga_row >= 10d"272" and vga_row < 10d"276") and (vga_col >= 10d"400" and vga_col < 10d"412")) or
								((vga_row >= 10d"276" and vga_row < 10d"280") and (vga_col >= 10d"232" and vga_col < 10d"244")) or
								((vga_row >= 10d"276" and vga_row < 10d"280") and (vga_col >= 10d"272" and vga_col < 10d"284")) or
								((vga_row >= 10d"276" and vga_row < 10d"280") and (vga_col >= 10d"300" and vga_col < 10d"312")) or
								((vga_row >= 10d"276" and vga_row < 10d"280") and (vga_col >= 10d"360" and vga_col < 10d"372")) or
								((vga_row >= 10d"276" and vga_row < 10d"280") and (vga_col >= 10d"404" and vga_col < 10d"416")) or
								((vga_row >= 10d"280" and vga_row < 10d"284") and (vga_col >= 10d"232" and vga_col < 10d"244")) or
								((vga_row >= 10d"280" and vga_row < 10d"284") and (vga_col >= 10d"268" and vga_col < 10d"284")) or
								((vga_row >= 10d"280" and vga_row < 10d"284") and (vga_col >= 10d"300" and vga_col < 10d"312")) or
								((vga_row >= 10d"280" and vga_row < 10d"284") and (vga_col >= 10d"360" and vga_col < 10d"372")) or
								((vga_row >= 10d"280" and vga_row < 10d"284") and (vga_col >= 10d"404" and vga_col < 10d"416")) or
								((vga_row >= 10d"284" and vga_row < 10d"288") and (vga_col >= 10d"232" and vga_col < 10d"280")) or
								((vga_row >= 10d"284" and vga_row < 10d"288") and (vga_col >= 10d"300" and vga_col < 10d"344")) or
								((vga_row >= 10d"284" and vga_row < 10d"288") and (vga_col >= 10d"360" and vga_col < 10d"372")) or
								((vga_row >= 10d"284" and vga_row < 10d"288") and (vga_col >= 10d"404" and vga_col < 10d"416")) or
								((vga_row >= 10d"288" and vga_row < 10d"292") and (vga_col >= 10d"232" and vga_col < 10d"276")) or
								((vga_row >= 10d"288" and vga_row < 10d"292") and (vga_col >= 10d"300" and vga_col < 10d"344")) or
								((vga_row >= 10d"288" and vga_row < 10d"292") and (vga_col >= 10d"360" and vga_col < 10d"372")) or
								((vga_row >= 10d"288" and vga_row < 10d"292") and (vga_col >= 10d"404" and vga_col < 10d"416")) or
								((vga_row >= 10d"292" and vga_row < 10d"296") and (vga_col >= 10d"232" and vga_col < 10d"268")) or
								((vga_row >= 10d"292" and vga_row < 10d"296") and (vga_col >= 10d"300" and vga_col < 10d"344")) or
								((vga_row >= 10d"292" and vga_row < 10d"296") and (vga_col >= 10d"360" and vga_col < 10d"372")) or
								((vga_row >= 10d"292" and vga_row < 10d"296") and (vga_col >= 10d"404" and vga_col < 10d"416")) or
								((vga_row >= 10d"296" and vga_row < 10d"300") and (vga_col >= 10d"232" and vga_col < 10d"244")) or
								((vga_row >= 10d"296" and vga_row < 10d"300") and (vga_col >= 10d"256" and vga_col < 10d"272")) or
								((vga_row >= 10d"296" and vga_row < 10d"300") and (vga_col >= 10d"300" and vga_col < 10d"312")) or
								((vga_row >= 10d"296" and vga_row < 10d"300") and (vga_col >= 10d"360" and vga_col < 10d"372")) or
								((vga_row >= 10d"296" and vga_row < 10d"300") and (vga_col >= 10d"404" and vga_col < 10d"416")) or
								((vga_row >= 10d"300" and vga_row < 10d"304") and (vga_col >= 10d"232" and vga_col < 10d"244")) or
								((vga_row >= 10d"300" and vga_row < 10d"304") and (vga_col >= 10d"260" and vga_col < 10d"276")) or
								((vga_row >= 10d"300" and vga_row < 10d"304") and (vga_col >= 10d"300" and vga_col < 10d"312")) or
								((vga_row >= 10d"300" and vga_row < 10d"304") and (vga_col >= 10d"360" and vga_col < 10d"372")) or
								((vga_row >= 10d"300" and vga_row < 10d"304") and (vga_col >= 10d"404" and vga_col < 10d"416")) or
								((vga_row >= 10d"304" and vga_row < 10d"308") and (vga_col >= 10d"232" and vga_col < 10d"244")) or
								((vga_row >= 10d"304" and vga_row < 10d"308") and (vga_col >= 10d"264" and vga_col < 10d"276")) or
								((vga_row >= 10d"304" and vga_row < 10d"308") and (vga_col >= 10d"300" and vga_col < 10d"312")) or
								((vga_row >= 10d"304" and vga_row < 10d"308") and (vga_col >= 10d"360" and vga_col < 10d"372")) or
								((vga_row >= 10d"304" and vga_row < 10d"308") and (vga_col >= 10d"400" and vga_col < 10d"412")) or
								((vga_row >= 10d"308" and vga_row < 10d"312") and (vga_col >= 10d"232" and vga_col < 10d"244")) or
								((vga_row >= 10d"308" and vga_row < 10d"312") and (vga_col >= 10d"268" and vga_col < 10d"280")) or
								((vga_row >= 10d"308" and vga_row < 10d"312") and (vga_col >= 10d"300" and vga_col < 10d"312")) or
								((vga_row >= 10d"308" and vga_row < 10d"312") and (vga_col >= 10d"360" and vga_col < 10d"372")) or
								((vga_row >= 10d"308" and vga_row < 10d"312") and (vga_col >= 10d"396" and vga_col < 10d"412")) or
								((vga_row >= 10d"312" and vga_row < 10d"316") and (vga_col >= 10d"232" and vga_col < 10d"244")) or
								((vga_row >= 10d"312" and vga_row < 10d"316") and (vga_col >= 10d"268" and vga_col < 10d"284")) or
								((vga_row >= 10d"312" and vga_row < 10d"316") and (vga_col >= 10d"300" and vga_col < 10d"348")) or
								((vga_row >= 10d"312" and vga_row < 10d"316") and (vga_col >= 10d"360" and vga_col < 10d"408")) or
								((vga_row >= 10d"316" and vga_row < 10d"320") and (vga_col >= 10d"232" and vga_col < 10d"244")) or
								((vga_row >= 10d"316" and vga_row < 10d"320") and (vga_col >= 10d"272" and vga_col < 10d"284")) or
								((vga_row >= 10d"316" and vga_row < 10d"320") and (vga_col >= 10d"300" and vga_col < 10d"348")) or
								((vga_row >= 10d"316" and vga_row < 10d"320") and (vga_col >= 10d"360" and vga_col < 10d"404")) or
								((vga_row >= 10d"320" and vga_row < 10d"324") and (vga_col >= 10d"232" and vga_col < 10d"244")) or
								((vga_row >= 10d"320" and vga_row < 10d"324") and (vga_col >= 10d"272" and vga_col < 10d"288")) or
								((vga_row >= 10d"320" and vga_row < 10d"324") and (vga_col >= 10d"300" and vga_col < 10d"348")) or
								((vga_row >= 10d"320" and vga_row < 10d"324") and (vga_col >= 10d"360" and vga_col < 10d"400"))) else
								
				 "000011" when player = '1' and 
								(((vga_row >= 10d"152" and vga_row < 10d"156") and (vga_col >= 10d"124" and vga_col < 10d"136")) or
								((vga_row >= 10d"152" and vga_row < 10d"156") and (vga_col >= 10d"160" and vga_col < 10d"172")) or
								((vga_row >= 10d"152" and vga_row < 10d"156") and (vga_col >= 10d"196" and vga_col < 10d"208")) or
								((vga_row >= 10d"152" and vga_row < 10d"156") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"152" and vga_row < 10d"156") and (vga_col >= 10d"236" and vga_col < 10d"248")) or
								((vga_row >= 10d"152" and vga_row < 10d"156") and (vga_col >= 10d"276" and vga_col < 10d"288")) or
								((vga_row >= 10d"152" and vga_row < 10d"156") and (vga_col >= 10d"304" and vga_col < 10d"316")) or
								((vga_row >= 10d"152" and vga_row < 10d"156") and (vga_col >= 10d"344" and vga_col < 10d"356")) or
								((vga_row >= 10d"152" and vga_row < 10d"156") and (vga_col >= 10d"372" and vga_col < 10d"420")) or
								((vga_row >= 10d"152" and vga_row < 10d"156") and (vga_col >= 10d"432" and vga_col < 10d"476")) or
								((vga_row >= 10d"156" and vga_row < 10d"160") and (vga_col >= 10d"124" and vga_col < 10d"136")) or
								((vga_row >= 10d"156" and vga_row < 10d"160") and (vga_col >= 10d"160" and vga_col < 10d"172")) or
								((vga_row >= 10d"156" and vga_row < 10d"160") and (vga_col >= 10d"196" and vga_col < 10d"208")) or
								((vga_row >= 10d"156" and vga_row < 10d"160") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"156" and vga_row < 10d"160") and (vga_col >= 10d"236" and vga_col < 10d"252")) or
								((vga_row >= 10d"156" and vga_row < 10d"160") and (vga_col >= 10d"276" and vga_col < 10d"288")) or
								((vga_row >= 10d"156" and vga_row < 10d"160") and (vga_col >= 10d"304" and vga_col < 10d"320")) or
								((vga_row >= 10d"156" and vga_row < 10d"160") and (vga_col >= 10d"344" and vga_col < 10d"356")) or
								((vga_row >= 10d"156" and vga_row < 10d"160") and (vga_col >= 10d"372" and vga_col < 10d"420")) or
								((vga_row >= 10d"156" and vga_row < 10d"160") and (vga_col >= 10d"432" and vga_col < 10d"480")) or
								((vga_row >= 10d"160" and vga_row < 10d"164") and (vga_col >= 10d"128" and vga_col < 10d"140")) or
								((vga_row >= 10d"160" and vga_row < 10d"164") and (vga_col >= 10d"156" and vga_col < 10d"176")) or
								((vga_row >= 10d"160" and vga_row < 10d"164") and (vga_col >= 10d"192" and vga_col < 10d"204")) or
								((vga_row >= 10d"160" and vga_row < 10d"164") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"160" and vga_row < 10d"164") and (vga_col >= 10d"236" and vga_col < 10d"256")) or
								((vga_row >= 10d"160" and vga_row < 10d"164") and (vga_col >= 10d"276" and vga_col < 10d"288")) or
								((vga_row >= 10d"160" and vga_row < 10d"164") and (vga_col >= 10d"304" and vga_col < 10d"324")) or
								((vga_row >= 10d"160" and vga_row < 10d"164") and (vga_col >= 10d"344" and vga_col < 10d"356")) or
								((vga_row >= 10d"160" and vga_row < 10d"164") and (vga_col >= 10d"372" and vga_col < 10d"420")) or
								((vga_row >= 10d"160" and vga_row < 10d"164") and (vga_col >= 10d"432" and vga_col < 10d"484")) or
								((vga_row >= 10d"164" and vga_row < 10d"168") and (vga_col >= 10d"128" and vga_col < 10d"140")) or
								((vga_row >= 10d"164" and vga_row < 10d"168") and (vga_col >= 10d"156" and vga_col < 10d"176")) or
								((vga_row >= 10d"164" and vga_row < 10d"168") and (vga_col >= 10d"192" and vga_col < 10d"204")) or
								((vga_row >= 10d"164" and vga_row < 10d"168") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"164" and vga_row < 10d"168") and (vga_col >= 10d"236" and vga_col < 10d"256")) or
								((vga_row >= 10d"164" and vga_row < 10d"168") and (vga_col >= 10d"276" and vga_col < 10d"288")) or
								((vga_row >= 10d"164" and vga_row < 10d"168") and (vga_col >= 10d"304" and vga_col < 10d"324")) or
								((vga_row >= 10d"164" and vga_row < 10d"168") and (vga_col >= 10d"344" and vga_col < 10d"356")) or
								((vga_row >= 10d"164" and vga_row < 10d"168") and (vga_col >= 10d"372" and vga_col < 10d"384")) or
								((vga_row >= 10d"164" and vga_row < 10d"168") and (vga_col >= 10d"432" and vga_col < 10d"444")) or
								((vga_row >= 10d"164" and vga_row < 10d"168") and (vga_col >= 10d"468" and vga_col < 10d"484")) or
								((vga_row >= 10d"168" and vga_row < 10d"172") and (vga_col >= 10d"128" and vga_col < 10d"140")) or
								((vga_row >= 10d"168" and vga_row < 10d"172") and (vga_col >= 10d"156" and vga_col < 10d"164")) or
								((vga_row >= 10d"168" and vga_row < 10d"172") and (vga_col >= 10d"168" and vga_col < 10d"176")) or
								((vga_row >= 10d"168" and vga_row < 10d"172") and (vga_col >= 10d"192" and vga_col < 10d"204")) or
								((vga_row >= 10d"168" and vga_row < 10d"172") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"168" and vga_row < 10d"172") and (vga_col >= 10d"236" and vga_col < 10d"260")) or
								((vga_row >= 10d"168" and vga_row < 10d"172") and (vga_col >= 10d"276" and vga_col < 10d"288")) or
								((vga_row >= 10d"168" and vga_row < 10d"172") and (vga_col >= 10d"304" and vga_col < 10d"328")) or
								((vga_row >= 10d"168" and vga_row < 10d"172") and (vga_col >= 10d"344" and vga_col < 10d"356")) or
								((vga_row >= 10d"168" and vga_row < 10d"172") and (vga_col >= 10d"372" and vga_col < 10d"384")) or
								((vga_row >= 10d"168" and vga_row < 10d"172") and (vga_col >= 10d"432" and vga_col < 10d"444")) or
								((vga_row >= 10d"168" and vga_row < 10d"172") and (vga_col >= 10d"472" and vga_col < 10d"484")) or
								((vga_row >= 10d"172" and vga_row < 10d"176") and (vga_col >= 10d"128" and vga_col < 10d"140")) or
								((vga_row >= 10d"172" and vga_row < 10d"176") and (vga_col >= 10d"152" and vga_col < 10d"164")) or
								((vga_row >= 10d"172" and vga_row < 10d"176") and (vga_col >= 10d"168" and vga_col < 10d"180")) or
								((vga_row >= 10d"172" and vga_row < 10d"176") and (vga_col >= 10d"192" and vga_col < 10d"204")) or
								((vga_row >= 10d"172" and vga_row < 10d"176") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"172" and vga_row < 10d"176") and (vga_col >= 10d"236" and vga_col < 10d"260")) or
								((vga_row >= 10d"172" and vga_row < 10d"176") and (vga_col >= 10d"276" and vga_col < 10d"288")) or
								((vga_row >= 10d"172" and vga_row < 10d"176") and (vga_col >= 10d"304" and vga_col < 10d"328")) or
								((vga_row >= 10d"172" and vga_row < 10d"176") and (vga_col >= 10d"344" and vga_col < 10d"356")) or
								((vga_row >= 10d"172" and vga_row < 10d"176") and (vga_col >= 10d"372" and vga_col < 10d"384")) or
								((vga_row >= 10d"172" and vga_row < 10d"176") and (vga_col >= 10d"432" and vga_col < 10d"444")) or
								((vga_row >= 10d"172" and vga_row < 10d"176") and (vga_col >= 10d"472" and vga_col < 10d"484")) or
								((vga_row >= 10d"172" and vga_row < 10d"176") and (vga_col >= 10d"500" and vga_col < 10d"512")) or
								((vga_row >= 10d"176" and vga_row < 10d"180") and (vga_col >= 10d"128" and vga_col < 10d"140")) or
								((vga_row >= 10d"176" and vga_row < 10d"180") and (vga_col >= 10d"152" and vga_col < 10d"164")) or
								((vga_row >= 10d"176" and vga_row < 10d"180") and (vga_col >= 10d"168" and vga_col < 10d"180")) or
								((vga_row >= 10d"176" and vga_row < 10d"180") and (vga_col >= 10d"192" and vga_col < 10d"204")) or
								((vga_row >= 10d"176" and vga_row < 10d"180") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"176" and vga_row < 10d"180") and (vga_col >= 10d"236" and vga_col < 10d"248")) or
								((vga_row >= 10d"176" and vga_row < 10d"180") and (vga_col >= 10d"252" and vga_col < 10d"264")) or
								((vga_row >= 10d"176" and vga_row < 10d"180") and (vga_col >= 10d"276" and vga_col < 10d"288")) or
								((vga_row >= 10d"176" and vga_row < 10d"180") and (vga_col >= 10d"304" and vga_col < 10d"316")) or
								((vga_row >= 10d"176" and vga_row < 10d"180") and (vga_col >= 10d"320" and vga_col < 10d"332")) or
								((vga_row >= 10d"176" and vga_row < 10d"180") and (vga_col >= 10d"344" and vga_col < 10d"356")) or
								((vga_row >= 10d"176" and vga_row < 10d"180") and (vga_col >= 10d"372" and vga_col < 10d"384")) or
								((vga_row >= 10d"176" and vga_row < 10d"180") and (vga_col >= 10d"432" and vga_col < 10d"444")) or
								((vga_row >= 10d"176" and vga_row < 10d"180") and (vga_col >= 10d"468" and vga_col < 10d"484")) or
								((vga_row >= 10d"176" and vga_row < 10d"180") and (vga_col >= 10d"500" and vga_col < 10d"512")) or
								((vga_row >= 10d"180" and vga_row < 10d"184") and (vga_col >= 10d"132" and vga_col < 10d"144")) or
								((vga_row >= 10d"180" and vga_row < 10d"184") and (vga_col >= 10d"152" and vga_col < 10d"164")) or
								((vga_row >= 10d"180" and vga_row < 10d"184") and (vga_col >= 10d"168" and vga_col < 10d"180")) or
								((vga_row >= 10d"180" and vga_row < 10d"184") and (vga_col >= 10d"188" and vga_col < 10d"200")) or
								((vga_row >= 10d"180" and vga_row < 10d"184") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"180" and vga_row < 10d"184") and (vga_col >= 10d"236" and vga_col < 10d"248")) or
								((vga_row >= 10d"180" and vga_row < 10d"184") and (vga_col >= 10d"252" and vga_col < 10d"264")) or
								((vga_row >= 10d"180" and vga_row < 10d"184") and (vga_col >= 10d"276" and vga_col < 10d"288")) or
								((vga_row >= 10d"180" and vga_row < 10d"184") and (vga_col >= 10d"304" and vga_col < 10d"316")) or
								((vga_row >= 10d"180" and vga_row < 10d"184") and (vga_col >= 10d"320" and vga_col < 10d"332")) or
								((vga_row >= 10d"180" and vga_row < 10d"184") and (vga_col >= 10d"344" and vga_col < 10d"356")) or
								((vga_row >= 10d"180" and vga_row < 10d"184") and (vga_col >= 10d"372" and vga_col < 10d"416")) or
								((vga_row >= 10d"180" and vga_row < 10d"184") and (vga_col >= 10d"432" and vga_col < 10d"480")) or
								((vga_row >= 10d"180" and vga_row < 10d"184") and (vga_col >= 10d"500" and vga_col < 10d"512")) or
								((vga_row >= 10d"184" and vga_row < 10d"188") and (vga_col >= 10d"132" and vga_col < 10d"144")) or
								((vga_row >= 10d"184" and vga_row < 10d"188") and (vga_col >= 10d"148" and vga_col < 10d"160")) or
								((vga_row >= 10d"184" and vga_row < 10d"188") and (vga_col >= 10d"172" and vga_col < 10d"180")) or
								((vga_row >= 10d"184" and vga_row < 10d"188") and (vga_col >= 10d"188" and vga_col < 10d"200")) or
								((vga_row >= 10d"184" and vga_row < 10d"188") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"184" and vga_row < 10d"188") and (vga_col >= 10d"236" and vga_col < 10d"248")) or
								((vga_row >= 10d"184" and vga_row < 10d"188") and (vga_col >= 10d"256" and vga_col < 10d"268")) or
								((vga_row >= 10d"184" and vga_row < 10d"188") and (vga_col >= 10d"276" and vga_col < 10d"288")) or
								((vga_row >= 10d"184" and vga_row < 10d"188") and (vga_col >= 10d"304" and vga_col < 10d"316")) or
								((vga_row >= 10d"184" and vga_row < 10d"188") and (vga_col >= 10d"324" and vga_col < 10d"336")) or
								((vga_row >= 10d"184" and vga_row < 10d"188") and (vga_col >= 10d"344" and vga_col < 10d"356")) or
								((vga_row >= 10d"184" and vga_row < 10d"188") and (vga_col >= 10d"372" and vga_col < 10d"416")) or
								((vga_row >= 10d"184" and vga_row < 10d"188") and (vga_col >= 10d"432" and vga_col < 10d"476")) or
								((vga_row >= 10d"188" and vga_row < 10d"192") and (vga_col >= 10d"132" and vga_col < 10d"144")) or
								((vga_row >= 10d"188" and vga_row < 10d"192") and (vga_col >= 10d"148" and vga_col < 10d"160")) or
								((vga_row >= 10d"188" and vga_row < 10d"192") and (vga_col >= 10d"172" and vga_col < 10d"184")) or
								((vga_row >= 10d"188" and vga_row < 10d"192") and (vga_col >= 10d"188" and vga_col < 10d"200")) or
								((vga_row >= 10d"188" and vga_row < 10d"192") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"188" and vga_row < 10d"192") and (vga_col >= 10d"236" and vga_col < 10d"248")) or
								((vga_row >= 10d"188" and vga_row < 10d"192") and (vga_col >= 10d"256" and vga_col < 10d"272")) or
								((vga_row >= 10d"188" and vga_row < 10d"192") and (vga_col >= 10d"276" and vga_col < 10d"288")) or
								((vga_row >= 10d"188" and vga_row < 10d"192") and (vga_col >= 10d"304" and vga_col < 10d"316")) or
								((vga_row >= 10d"188" and vga_row < 10d"192") and (vga_col >= 10d"324" and vga_col < 10d"340")) or
								((vga_row >= 10d"188" and vga_row < 10d"192") and (vga_col >= 10d"344" and vga_col < 10d"356")) or
								((vga_row >= 10d"188" and vga_row < 10d"192") and (vga_col >= 10d"372" and vga_col < 10d"416")) or
								((vga_row >= 10d"188" and vga_row < 10d"192") and (vga_col >= 10d"432" and vga_col < 10d"468")) or
								((vga_row >= 10d"192" and vga_row < 10d"196") and (vga_col >= 10d"132" and vga_col < 10d"144")) or
								((vga_row >= 10d"192" and vga_row < 10d"196") and (vga_col >= 10d"148" and vga_col < 10d"160")) or
								((vga_row >= 10d"192" and vga_row < 10d"196") and (vga_col >= 10d"172" and vga_col < 10d"184")) or
								((vga_row >= 10d"192" and vga_row < 10d"196") and (vga_col >= 10d"188" and vga_col < 10d"200")) or
								((vga_row >= 10d"192" and vga_row < 10d"196") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"192" and vga_row < 10d"196") and (vga_col >= 10d"236" and vga_col < 10d"248")) or
								((vga_row >= 10d"192" and vga_row < 10d"196") and (vga_col >= 10d"260" and vga_col < 10d"272")) or
								((vga_row >= 10d"192" and vga_row < 10d"196") and (vga_col >= 10d"276" and vga_col < 10d"288")) or
								((vga_row >= 10d"192" and vga_row < 10d"196") and (vga_col >= 10d"304" and vga_col < 10d"316")) or
								((vga_row >= 10d"192" and vga_row < 10d"196") and (vga_col >= 10d"328" and vga_col < 10d"340")) or
								((vga_row >= 10d"192" and vga_row < 10d"196") and (vga_col >= 10d"344" and vga_col < 10d"356")) or
								((vga_row >= 10d"192" and vga_row < 10d"196") and (vga_col >= 10d"372" and vga_col < 10d"384")) or
								((vga_row >= 10d"192" and vga_row < 10d"196") and (vga_col >= 10d"432" and vga_col < 10d"444")) or
								((vga_row >= 10d"192" and vga_row < 10d"196") and (vga_col >= 10d"456" and vga_col < 10d"472")) or
								((vga_row >= 10d"196" and vga_row < 10d"200") and (vga_col >= 10d"136" and vga_col < 10d"144")) or
								((vga_row >= 10d"196" and vga_row < 10d"200") and (vga_col >= 10d"148" and vga_col < 10d"160")) or
								((vga_row >= 10d"196" and vga_row < 10d"200") and (vga_col >= 10d"172" and vga_col < 10d"184")) or
								((vga_row >= 10d"196" and vga_row < 10d"200") and (vga_col >= 10d"188" and vga_col < 10d"196")) or
								((vga_row >= 10d"196" and vga_row < 10d"200") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"196" and vga_row < 10d"200") and (vga_col >= 10d"236" and vga_col < 10d"248")) or
								((vga_row >= 10d"196" and vga_row < 10d"200") and (vga_col >= 10d"264" and vga_col < 10d"288")) or
								((vga_row >= 10d"196" and vga_row < 10d"200") and (vga_col >= 10d"304" and vga_col < 10d"316")) or
								((vga_row >= 10d"196" and vga_row < 10d"200") and (vga_col >= 10d"332" and vga_col < 10d"356")) or
								((vga_row >= 10d"196" and vga_row < 10d"200") and (vga_col >= 10d"372" and vga_col < 10d"384")) or
								((vga_row >= 10d"196" and vga_row < 10d"200") and (vga_col >= 10d"432" and vga_col < 10d"444")) or
								((vga_row >= 10d"196" and vga_row < 10d"200") and (vga_col >= 10d"460" and vga_col < 10d"476")) or
								((vga_row >= 10d"200" and vga_row < 10d"204") and (vga_col >= 10d"136" and vga_col < 10d"156")) or
								((vga_row >= 10d"200" and vga_row < 10d"204") and (vga_col >= 10d"176" and vga_col < 10d"196")) or
								((vga_row >= 10d"200" and vga_row < 10d"204") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"200" and vga_row < 10d"204") and (vga_col >= 10d"236" and vga_col < 10d"248")) or
								((vga_row >= 10d"200" and vga_row < 10d"204") and (vga_col >= 10d"264" and vga_col < 10d"288")) or
								((vga_row >= 10d"200" and vga_row < 10d"204") and (vga_col >= 10d"304" and vga_col < 10d"316")) or
								((vga_row >= 10d"200" and vga_row < 10d"204") and (vga_col >= 10d"332" and vga_col < 10d"356")) or
								((vga_row >= 10d"200" and vga_row < 10d"204") and (vga_col >= 10d"372" and vga_col < 10d"384")) or
								((vga_row >= 10d"200" and vga_row < 10d"204") and (vga_col >= 10d"432" and vga_col < 10d"444")) or
								((vga_row >= 10d"200" and vga_row < 10d"204") and (vga_col >= 10d"464" and vga_col < 10d"476")) or
								((vga_row >= 10d"204" and vga_row < 10d"208") and (vga_col >= 10d"136" and vga_col < 10d"156")) or
								((vga_row >= 10d"204" and vga_row < 10d"208") and (vga_col >= 10d"176" and vga_col < 10d"196")) or
								((vga_row >= 10d"204" and vga_row < 10d"208") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"204" and vga_row < 10d"208") and (vga_col >= 10d"236" and vga_col < 10d"248")) or
								((vga_row >= 10d"204" and vga_row < 10d"208") and (vga_col >= 10d"268" and vga_col < 10d"288")) or
								((vga_row >= 10d"204" and vga_row < 10d"208") and (vga_col >= 10d"304" and vga_col < 10d"316")) or
								((vga_row >= 10d"204" and vga_row < 10d"208") and (vga_col >= 10d"336" and vga_col < 10d"356")) or
								((vga_row >= 10d"204" and vga_row < 10d"208") and (vga_col >= 10d"372" and vga_col < 10d"384")) or
								((vga_row >= 10d"204" and vga_row < 10d"208") and (vga_col >= 10d"432" and vga_col < 10d"444")) or
								((vga_row >= 10d"204" and vga_row < 10d"208") and (vga_col >= 10d"468" and vga_col < 10d"480")) or
								((vga_row >= 10d"208" and vga_row < 10d"212") and (vga_col >= 10d"136" and vga_col < 10d"156")) or
								((vga_row >= 10d"208" and vga_row < 10d"212") and (vga_col >= 10d"176" and vga_col < 10d"196")) or
								((vga_row >= 10d"208" and vga_row < 10d"212") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"208" and vga_row < 10d"212") and (vga_col >= 10d"236" and vga_col < 10d"248")) or
								((vga_row >= 10d"208" and vga_row < 10d"212") and (vga_col >= 10d"268" and vga_col < 10d"288")) or
								((vga_row >= 10d"208" and vga_row < 10d"212") and (vga_col >= 10d"304" and vga_col < 10d"316")) or
								((vga_row >= 10d"208" and vga_row < 10d"212") and (vga_col >= 10d"336" and vga_col < 10d"356")) or
								((vga_row >= 10d"208" and vga_row < 10d"212") and (vga_col >= 10d"372" and vga_col < 10d"420")) or
								((vga_row >= 10d"208" and vga_row < 10d"212") and (vga_col >= 10d"432" and vga_col < 10d"444")) or
								((vga_row >= 10d"208" and vga_row < 10d"212") and (vga_col >= 10d"468" and vga_col < 10d"484")) or
								((vga_row >= 10d"208" and vga_row < 10d"212") and (vga_col >= 10d"500" and vga_col < 10d"512")) or
								((vga_row >= 10d"212" and vga_row < 10d"216") and (vga_col >= 10d"140" and vga_col < 10d"152")) or
								((vga_row >= 10d"212" and vga_row < 10d"216") and (vga_col >= 10d"180" and vga_col < 10d"192")) or
								((vga_row >= 10d"212" and vga_row < 10d"216") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"212" and vga_row < 10d"216") and (vga_col >= 10d"236" and vga_col < 10d"248")) or
								((vga_row >= 10d"212" and vga_row < 10d"216") and (vga_col >= 10d"272" and vga_col < 10d"288")) or
								((vga_row >= 10d"212" and vga_row < 10d"216") and (vga_col >= 10d"304" and vga_col < 10d"316")) or
								((vga_row >= 10d"212" and vga_row < 10d"216") and (vga_col >= 10d"340" and vga_col < 10d"356")) or
								((vga_row >= 10d"212" and vga_row < 10d"216") and (vga_col >= 10d"372" and vga_col < 10d"420")) or
								((vga_row >= 10d"212" and vga_row < 10d"216") and (vga_col >= 10d"432" and vga_col < 10d"444")) or
								((vga_row >= 10d"212" and vga_row < 10d"216") and (vga_col >= 10d"472" and vga_col < 10d"484")) or
								((vga_row >= 10d"212" and vga_row < 10d"216") and (vga_col >= 10d"500" and vga_col < 10d"512")) or
								((vga_row >= 10d"216" and vga_row < 10d"220") and (vga_col >= 10d"140" and vga_col < 10d"152")) or
								((vga_row >= 10d"216" and vga_row < 10d"220") and (vga_col >= 10d"180" and vga_col < 10d"192")) or
								((vga_row >= 10d"216" and vga_row < 10d"220") and (vga_col >= 10d"212" and vga_col < 10d"224")) or
								((vga_row >= 10d"216" and vga_row < 10d"220") and (vga_col >= 10d"236" and vga_col < 10d"248")) or
								((vga_row >= 10d"216" and vga_row < 10d"220") and (vga_col >= 10d"272" and vga_col < 10d"288")) or
								((vga_row >= 10d"216" and vga_row < 10d"220") and (vga_col >= 10d"304" and vga_col < 10d"316")) or
								((vga_row >= 10d"216" and vga_row < 10d"220") and (vga_col >= 10d"340" and vga_col < 10d"356")) or
								((vga_row >= 10d"216" and vga_row < 10d"220") and (vga_col >= 10d"372" and vga_col < 10d"420")) or
								((vga_row >= 10d"216" and vga_row < 10d"220") and (vga_col >= 10d"432" and vga_col < 10d"444")) or
								((vga_row >= 10d"216" and vga_row < 10d"220") and (vga_col >= 10d"472" and vga_col < 10d"488")) or
								((vga_row >= 10d"216" and vga_row < 10d"220") and (vga_col >= 10d"500" and vga_col < 10d"512")) or
								((vga_row >= 10d"256" and vga_row < 10d"260") and (vga_col >= 10d"204" and vga_col < 10d"248")) or
								((vga_row >= 10d"256" and vga_row < 10d"260") and (vga_col >= 10d"272" and vga_col < 10d"284")) or
								((vga_row >= 10d"256" and vga_row < 10d"260") and (vga_col >= 10d"328" and vga_col < 10d"340")) or
								((vga_row >= 10d"256" and vga_row < 10d"260") and (vga_col >= 10d"368" and vga_col < 10d"380")) or
								((vga_row >= 10d"256" and vga_row < 10d"260") and (vga_col >= 10d"396" and vga_col < 10d"444")) or
								((vga_row >= 10d"260" and vga_row < 10d"264") and (vga_col >= 10d"204" and vga_col < 10d"252")) or
								((vga_row >= 10d"260" and vga_row < 10d"264") and (vga_col >= 10d"272" and vga_col < 10d"284")) or
								((vga_row >= 10d"260" and vga_row < 10d"264") and (vga_col >= 10d"328" and vga_col < 10d"340")) or
								((vga_row >= 10d"260" and vga_row < 10d"264") and (vga_col >= 10d"368" and vga_col < 10d"380")) or
								((vga_row >= 10d"260" and vga_row < 10d"264") and (vga_col >= 10d"396" and vga_col < 10d"444")) or
								((vga_row >= 10d"264" and vga_row < 10d"268") and (vga_col >= 10d"204" and vga_col < 10d"252")) or
								((vga_row >= 10d"264" and vga_row < 10d"268") and (vga_col >= 10d"272" and vga_col < 10d"284")) or
								((vga_row >= 10d"264" and vga_row < 10d"268") and (vga_col >= 10d"328" and vga_col < 10d"340")) or
								((vga_row >= 10d"264" and vga_row < 10d"268") and (vga_col >= 10d"368" and vga_col < 10d"380")) or
								((vga_row >= 10d"264" and vga_row < 10d"268") and (vga_col >= 10d"396" and vga_col < 10d"444")) or
								((vga_row >= 10d"268" and vga_row < 10d"272") and (vga_col >= 10d"204" and vga_col < 10d"216")) or
								((vga_row >= 10d"268" and vga_row < 10d"272") and (vga_col >= 10d"240" and vga_col < 10d"256")) or
								((vga_row >= 10d"268" and vga_row < 10d"272") and (vga_col >= 10d"272" and vga_col < 10d"284")) or
								((vga_row >= 10d"268" and vga_row < 10d"272") and (vga_col >= 10d"328" and vga_col < 10d"340")) or
								((vga_row >= 10d"268" and vga_row < 10d"272") and (vga_col >= 10d"368" and vga_col < 10d"380")) or
								((vga_row >= 10d"268" and vga_row < 10d"272") and (vga_col >= 10d"396" and vga_col < 10d"408")) or
								((vga_row >= 10d"272" and vga_row < 10d"276") and (vga_col >= 10d"204" and vga_col < 10d"216")) or
								((vga_row >= 10d"272" and vga_row < 10d"276") and (vga_col >= 10d"244" and vga_col < 10d"256")) or
								((vga_row >= 10d"272" and vga_row < 10d"276") and (vga_col >= 10d"272" and vga_col < 10d"284")) or
								((vga_row >= 10d"272" and vga_row < 10d"276") and (vga_col >= 10d"328" and vga_col < 10d"340")) or
								((vga_row >= 10d"272" and vga_row < 10d"276") and (vga_col >= 10d"368" and vga_col < 10d"380")) or
								((vga_row >= 10d"272" and vga_row < 10d"276") and (vga_col >= 10d"396" and vga_col < 10d"408")) or
								((vga_row >= 10d"276" and vga_row < 10d"280") and (vga_col >= 10d"204" and vga_col < 10d"216")) or
								((vga_row >= 10d"276" and vga_row < 10d"280") and (vga_col >= 10d"244" and vga_col < 10d"256")) or
								((vga_row >= 10d"276" and vga_row < 10d"280") and (vga_col >= 10d"272" and vga_col < 10d"284")) or
								((vga_row >= 10d"276" and vga_row < 10d"280") and (vga_col >= 10d"328" and vga_col < 10d"340")) or
								((vga_row >= 10d"276" and vga_row < 10d"280") and (vga_col >= 10d"368" and vga_col < 10d"380")) or
								((vga_row >= 10d"276" and vga_row < 10d"280") and (vga_col >= 10d"396" and vga_col < 10d"408")) or
								((vga_row >= 10d"280" and vga_row < 10d"284") and (vga_col >= 10d"204" and vga_col < 10d"216")) or
								((vga_row >= 10d"280" and vga_row < 10d"284") and (vga_col >= 10d"240" and vga_col < 10d"256")) or
								((vga_row >= 10d"280" and vga_row < 10d"284") and (vga_col >= 10d"272" and vga_col < 10d"284")) or
								((vga_row >= 10d"280" and vga_row < 10d"284") and (vga_col >= 10d"328" and vga_col < 10d"340")) or
								((vga_row >= 10d"280" and vga_row < 10d"284") and (vga_col >= 10d"368" and vga_col < 10d"380")) or
								((vga_row >= 10d"280" and vga_row < 10d"284") and (vga_col >= 10d"396" and vga_col < 10d"408")) or
								((vga_row >= 10d"284" and vga_row < 10d"288") and (vga_col >= 10d"204" and vga_col < 10d"252")) or
								((vga_row >= 10d"284" and vga_row < 10d"288") and (vga_col >= 10d"272" and vga_col < 10d"284")) or
								((vga_row >= 10d"284" and vga_row < 10d"288") and (vga_col >= 10d"328" and vga_col < 10d"340")) or
								((vga_row >= 10d"284" and vga_row < 10d"288") and (vga_col >= 10d"368" and vga_col < 10d"380")) or
								((vga_row >= 10d"284" and vga_row < 10d"288") and (vga_col >= 10d"396" and vga_col < 10d"440")) or
								((vga_row >= 10d"288" and vga_row < 10d"292") and (vga_col >= 10d"204" and vga_col < 10d"252")) or
								((vga_row >= 10d"288" and vga_row < 10d"292") and (vga_col >= 10d"272" and vga_col < 10d"284")) or
								((vga_row >= 10d"288" and vga_row < 10d"292") and (vga_col >= 10d"328" and vga_col < 10d"340")) or
								((vga_row >= 10d"288" and vga_row < 10d"292") and (vga_col >= 10d"368" and vga_col < 10d"380")) or
								((vga_row >= 10d"288" and vga_row < 10d"292") and (vga_col >= 10d"396" and vga_col < 10d"440")) or
								((vga_row >= 10d"292" and vga_row < 10d"296") and (vga_col >= 10d"204" and vga_col < 10d"256")) or
								((vga_row >= 10d"292" and vga_row < 10d"296") and (vga_col >= 10d"272" and vga_col < 10d"284")) or
								((vga_row >= 10d"292" and vga_row < 10d"296") and (vga_col >= 10d"328" and vga_col < 10d"340")) or
								((vga_row >= 10d"292" and vga_row < 10d"296") and (vga_col >= 10d"368" and vga_col < 10d"380")) or
								((vga_row >= 10d"292" and vga_row < 10d"296") and (vga_col >= 10d"396" and vga_col < 10d"440")) or
								((vga_row >= 10d"296" and vga_row < 10d"300") and (vga_col >= 10d"204" and vga_col < 10d"216")) or
								((vga_row >= 10d"296" and vga_row < 10d"300") and (vga_col >= 10d"244" and vga_col < 10d"260")) or
								((vga_row >= 10d"296" and vga_row < 10d"300") and (vga_col >= 10d"272" and vga_col < 10d"284")) or
								((vga_row >= 10d"296" and vga_row < 10d"300") and (vga_col >= 10d"328" and vga_col < 10d"340")) or
								((vga_row >= 10d"296" and vga_row < 10d"300") and (vga_col >= 10d"368" and vga_col < 10d"380")) or
								((vga_row >= 10d"296" and vga_row < 10d"300") and (vga_col >= 10d"396" and vga_col < 10d"408")) or
								((vga_row >= 10d"300" and vga_row < 10d"304") and (vga_col >= 10d"204" and vga_col < 10d"216")) or
								((vga_row >= 10d"300" and vga_row < 10d"304") and (vga_col >= 10d"248" and vga_col < 10d"260")) or
								((vga_row >= 10d"300" and vga_row < 10d"304") and (vga_col >= 10d"272" and vga_col < 10d"284")) or
								((vga_row >= 10d"300" and vga_row < 10d"304") and (vga_col >= 10d"328" and vga_col < 10d"340")) or
								((vga_row >= 10d"300" and vga_row < 10d"304") and (vga_col >= 10d"368" and vga_col < 10d"380")) or
								((vga_row >= 10d"300" and vga_row < 10d"304") and (vga_col >= 10d"396" and vga_col < 10d"408")) or
								((vga_row >= 10d"304" and vga_row < 10d"308") and (vga_col >= 10d"204" and vga_col < 10d"216")) or
								((vga_row >= 10d"304" and vga_row < 10d"308") and (vga_col >= 10d"248" and vga_col < 10d"260")) or
								((vga_row >= 10d"304" and vga_row < 10d"308") and (vga_col >= 10d"272" and vga_col < 10d"284")) or
								((vga_row >= 10d"304" and vga_row < 10d"308") and (vga_col >= 10d"328" and vga_col < 10d"340")) or
								((vga_row >= 10d"304" and vga_row < 10d"308") and (vga_col >= 10d"368" and vga_col < 10d"380")) or
								((vga_row >= 10d"304" and vga_row < 10d"308") and (vga_col >= 10d"396" and vga_col < 10d"408")) or
								((vga_row >= 10d"308" and vga_row < 10d"312") and (vga_col >= 10d"204" and vga_col < 10d"216")) or
								((vga_row >= 10d"308" and vga_row < 10d"312") and (vga_col >= 10d"244" and vga_col < 10d"260")) or
								((vga_row >= 10d"308" and vga_row < 10d"312") and (vga_col >= 10d"272" and vga_col < 10d"284")) or
								((vga_row >= 10d"308" and vga_row < 10d"312") and (vga_col >= 10d"328" and vga_col < 10d"344")) or
								((vga_row >= 10d"308" and vga_row < 10d"312") and (vga_col >= 10d"364" and vga_col < 10d"380")) or
								((vga_row >= 10d"308" and vga_row < 10d"312") and (vga_col >= 10d"396" and vga_col < 10d"408")) or
								((vga_row >= 10d"312" and vga_row < 10d"316") and (vga_col >= 10d"204" and vga_col < 10d"256")) or
								((vga_row >= 10d"312" and vga_row < 10d"316") and (vga_col >= 10d"272" and vga_col < 10d"316")) or
								((vga_row >= 10d"312" and vga_row < 10d"316") and (vga_col >= 10d"332" and vga_col < 10d"376")) or
								((vga_row >= 10d"312" and vga_row < 10d"316") and (vga_col >= 10d"396" and vga_col < 10d"444")) or
								((vga_row >= 10d"316" and vga_row < 10d"320") and (vga_col >= 10d"204" and vga_col < 10d"256")) or
								((vga_row >= 10d"316" and vga_row < 10d"320") and (vga_col >= 10d"272" and vga_col < 10d"316")) or
								((vga_row >= 10d"316" and vga_row < 10d"320") and (vga_col >= 10d"336" and vga_col < 10d"372")) or
								((vga_row >= 10d"316" and vga_row < 10d"320") and (vga_col >= 10d"396" and vga_col < 10d"444")) or
								((vga_row >= 10d"320" and vga_row < 10d"324") and (vga_col >= 10d"204" and vga_col < 10d"248")) or
								((vga_row >= 10d"320" and vga_row < 10d"324") and (vga_col >= 10d"272" and vga_col < 10d"316")) or
								((vga_row >= 10d"320" and vga_row < 10d"324") and (vga_col >= 10d"340" and vga_col < 10d"368")) or
								((vga_row >= 10d"320" and vga_row < 10d"324") and (vga_col >= 10d"396" and vga_col < 10d"444"))) else
								"000000";
								
end;
